-- Elementos de Sistemas
-- by Rafael Corsi
-- MultiplicadorAcomB.vhd

Library ieee;
use ieee.std_logic_1164.all;

entity MultiplicadorAcomB is
	port(
		A     : in  STD_LOGIC_VECTOR(15 downto 0);
		B     : in  STD_LOGIC_VECTOR(15 downto 0);
		Y     : out STD_LOGIC_VECTOR(15 downto 0)
	);
end entity;

architecture arch of MultiplicadorAcomB is

begin

end architecture;
